LIBRARY IEEE;
USE IEEE.Std_Logic_1164.ALL;

ENTITY aritmetico IS
	PORT (
		A : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		B : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		SEL : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		OUTHEX : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		OUTBIN : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END aritmetico;

ARCHITECTURE arch OF aritmetico IS
	SIGNAL F1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL F2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL F3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL F4 : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL FMUX : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL G : STD_LOGIC_VECTOR(3 DOWNTO 0);
	COMPONENT somador IS
		PORT (
			A : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			F : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT mux IS
		PORT (
			W : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			X : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			Y : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			Z : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			SEL : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			F : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT decod7seg IS
		PORT (
			INPUT : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			HEX0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT circuito1 IS
		PORT (
			A : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			B : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			F1 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			F2 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			F3 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			F4 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
		);
	END COMPONENT;
BEGIN
	C1 : circuito1 PORT MAP(A, B, F1, F2, F3, F4);
	CMUX : mux PORT MAP(F1, F2, F3, F4, SEL, FMUX);
	CSUM : somador PORT MAP(F1, FMUX, G);
	CHEX : decod7seg PORT MAP(G, OUTHEX);
	OUTBIN <= G;
END arch;

